<?xml version='1.0' encoding='UTF-8'?> 
            <!DOCTYPE svg PUBLIC '-//W3C//DTD SVG 1.1//EN' 
            'http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd'>
<svg width='7505' height='3299' 
            xmlns='http://www.w3.org/2000/svg' version='1.1'>
<g><g style='font-family: "Sans";'>
<g transform='translate(10.000000, 0.000000) ' >
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3640.000000,2196.500000 4340.000000,2109.000000 4340.000000,2189.000000 3640.000000,2276.500000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1240.000000,2782.437500 1540.000000,2559.000000 1540.000000,2639.000000 1240.000000,2862.437500 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='640.000000,883.926758 840.000000,1708.853516 840.000000,1788.853516 640.000000,963.926758 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='0.000000,883.926758 640.000000,883.926758 640.000000,963.926758 0.000000,963.926758 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='640.000000,883.926758 740.000000,59.000000 740.000000,139.000000 640.000000,963.926758 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='5240.000000,2359.000000 6140.000000,2309.000000 6140.000000,2389.000000 5240.000000,2439.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1440.000000,1011.539062 2040.000000,1539.078125 2040.000000,1619.078125 1440.000000,1091.539062 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1440.000000,1011.539062 1940.000000,484.000000 1940.000000,564.000000 1440.000000,1091.539062 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='6340.000000,1059.000000 6540.000000,1009.000000 6540.000000,1089.000000 6340.000000,1139.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3840.000000,2984.000000 4640.000000,3059.000000 4640.000000,3139.000000 3840.000000,3064.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1140.000000,635.269531 1440.000000,1011.539062 1440.000000,1091.539062 1140.000000,715.269531 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1140.000000,635.269531 1340.000000,259.000000 1340.000000,339.000000 1140.000000,715.269531 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='840.000000,1708.853516 1240.000000,2782.437500 1240.000000,2862.437500 840.000000,1788.853516 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='840.000000,1708.853516 1140.000000,635.269531 1140.000000,715.269531 840.000000,1788.853516 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4440.000000,2284.000000 5240.000000,2359.000000 5240.000000,2439.000000 4440.000000,2364.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3840.000000,2984.000000 4540.000000,2909.000000 4540.000000,2989.000000 3840.000000,3064.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='740.000000,59.000000 940.000000,9.000000 940.000000,89.000000 740.000000,139.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1340.000000,259.000000 1840.000000,309.000000 1840.000000,389.000000 1340.000000,339.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2640.000000,559.000000 3140.000000,509.000000 3140.000000,589.000000 2640.000000,639.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4940.000000,1559.000000 5740.000000,1509.000000 5740.000000,1589.000000 4940.000000,1639.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4440.000000,2284.000000 5140.000000,2209.000000 5140.000000,2289.000000 4440.000000,2364.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1940.000000,484.000000 2540.000000,409.000000 2540.000000,489.000000 1940.000000,564.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='6440.000000,1284.000000 6840.000000,1359.000000 6840.000000,1439.000000 6440.000000,1364.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3540.000000,1959.000000 4240.000000,2009.000000 4240.000000,2089.000000 3540.000000,2039.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3640.000000,2196.500000 4440.000000,2284.000000 4440.000000,2364.000000 3640.000000,2276.500000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2740.000000,1000.406250 3440.000000,1291.812500 3440.000000,1371.812500 2740.000000,1080.406250 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='5640.000000,1171.500000 6340.000000,1059.000000 6340.000000,1139.000000 5640.000000,1251.500000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1640.000000,3005.875000 2340.000000,2802.750000 2340.000000,2882.750000 1640.000000,3085.875000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='5640.000000,1171.500000 6440.000000,1284.000000 6440.000000,1364.000000 5640.000000,1251.500000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3440.000000,1291.812500 4040.000000,1659.000000 4040.000000,1739.000000 3440.000000,1371.812500 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3440.000000,1291.812500 3940.000000,924.625000 3940.000000,1004.625000 3440.000000,1371.812500 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='6440.000000,1284.000000 6740.000000,1209.000000 6740.000000,1289.000000 6440.000000,1364.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3940.000000,924.625000 4740.000000,809.000000 4740.000000,889.000000 3940.000000,1004.625000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2640.000000,559.000000 3240.000000,609.000000 3240.000000,689.000000 2640.000000,639.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4640.000000,3059.000000 5440.000000,3109.000000 5440.000000,3189.000000 4640.000000,3139.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4840.000000,1040.250000 5540.000000,909.000000 5540.000000,989.000000 4840.000000,1120.250000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3540.000000,1959.000000 4140.000000,1909.000000 4140.000000,1989.000000 3540.000000,2039.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2340.000000,2802.750000 2940.000000,2709.000000 2940.000000,2789.000000 2340.000000,2882.750000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='740.000000,59.000000 1040.000000,109.000000 1040.000000,189.000000 740.000000,139.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1540.000000,2559.000000 2240.000000,2609.000000 2240.000000,2689.000000 1540.000000,2639.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2740.000000,1000.406250 3340.000000,709.000000 3340.000000,789.000000 2740.000000,1080.406250 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='5240.000000,2359.000000 6240.000000,2409.000000 6240.000000,2489.000000 5240.000000,2439.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4940.000000,1559.000000 5840.000000,1609.000000 5840.000000,1689.000000 4940.000000,1639.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1240.000000,2782.437500 1640.000000,3005.875000 1640.000000,3085.875000 1240.000000,2862.437500 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2840.000000,2077.750000 3540.000000,1959.000000 3540.000000,2039.000000 2840.000000,2157.750000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2840.000000,2077.750000 3640.000000,2196.500000 3640.000000,2276.500000 2840.000000,2157.750000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2040.000000,1539.078125 2740.000000,1000.406250 2740.000000,1080.406250 2040.000000,1619.078125 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2040.000000,1539.078125 2840.000000,2077.750000 2840.000000,2157.750000 2040.000000,1619.078125 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3040.000000,2896.500000 3840.000000,2984.000000 3840.000000,3064.000000 3040.000000,2976.500000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1940.000000,484.000000 2640.000000,559.000000 2640.000000,639.000000 1940.000000,564.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1540.000000,2559.000000 2140.000000,2509.000000 2140.000000,2589.000000 1540.000000,2639.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='6840.000000,1359.000000 7040.000000,1409.000000 7040.000000,1489.000000 6840.000000,1439.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1340.000000,259.000000 1740.000000,209.000000 1740.000000,289.000000 1340.000000,339.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='5040.000000,1759.000000 6040.000000,1809.000000 6040.000000,1889.000000 5040.000000,1839.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='1640.000000,3005.875000 2440.000000,3209.000000 2440.000000,3289.000000 1640.000000,3085.875000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3040.000000,2896.500000 3740.000000,2809.000000 3740.000000,2889.000000 3040.000000,2976.500000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4040.000000,1659.000000 4940.000000,1559.000000 4940.000000,1639.000000 4040.000000,1739.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4040.000000,1659.000000 5040.000000,1759.000000 5040.000000,1839.000000 4040.000000,1739.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='6340.000000,1059.000000 6640.000000,1109.000000 6640.000000,1189.000000 6340.000000,1139.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='2340.000000,2802.750000 3040.000000,2896.500000 3040.000000,2976.500000 2340.000000,2882.750000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='5040.000000,1759.000000 5940.000000,1709.000000 5940.000000,1789.000000 5040.000000,1839.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='3940.000000,924.625000 4840.000000,1040.250000 4840.000000,1120.250000 3940.000000,1004.625000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4840.000000,1040.250000 5640.000000,1171.500000 5640.000000,1251.500000 4840.000000,1120.250000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='6840.000000,1359.000000 6940.000000,1309.000000 6940.000000,1389.000000 6840.000000,1439.000000 ' stroke-width='1.000000'/>
<polygon stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(76,178,76)'  points='4640.000000,3059.000000 5340.000000,3009.000000 5340.000000,3089.000000 4640.000000,3139.000000 ' stroke-width='1.000000'/>
<line x1='1540.000000' y1='2559.000000' x2='1540.000000' y2='2639.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='840.000000' y1='1708.853516' x2='840.000000' y2='1788.853516' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='640.000000' y1='883.926758' x2='640.000000' y2='963.926758' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='740.000000' y1='59.000000' x2='740.000000' y2='139.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='2040.000000' y1='1539.078125' x2='2040.000000' y2='1619.078125' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='1940.000000' y1='484.000000' x2='1940.000000' y2='564.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='4640.000000' y1='3059.000000' x2='4640.000000' y2='3139.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='1440.000000' y1='1011.539062' x2='1440.000000' y2='1091.539062' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='1340.000000' y1='259.000000' x2='1340.000000' y2='339.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='1240.000000' y1='2782.437500' x2='1240.000000' y2='2862.437500' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='1140.000000' y1='635.269531' x2='1140.000000' y2='715.269531' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='5240.000000' y1='2359.000000' x2='5240.000000' y2='2439.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='6840.000000' y1='1359.000000' x2='6840.000000' y2='1439.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='4440.000000' y1='2284.000000' x2='4440.000000' y2='2364.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='3440.000000' y1='1291.812500' x2='3440.000000' y2='1371.812500' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='6340.000000' y1='1059.000000' x2='6340.000000' y2='1139.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='2340.000000' y1='2802.750000' x2='2340.000000' y2='2882.750000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='6440.000000' y1='1284.000000' x2='6440.000000' y2='1364.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='4040.000000' y1='1659.000000' x2='4040.000000' y2='1739.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='3940.000000' y1='924.625000' x2='3940.000000' y2='1004.625000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='1640.000000' y1='3005.875000' x2='1640.000000' y2='3085.875000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='3540.000000' y1='1959.000000' x2='3540.000000' y2='2039.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='3640.000000' y1='2196.500000' x2='3640.000000' y2='2276.500000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='2740.000000' y1='1000.406250' x2='2740.000000' y2='1080.406250' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='2840.000000' y1='2077.750000' x2='2840.000000' y2='2157.750000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='3840.000000' y1='2984.000000' x2='3840.000000' y2='3064.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='2640.000000' y1='559.000000' x2='2640.000000' y2='639.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='4940.000000' y1='1559.000000' x2='4940.000000' y2='1639.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='5040.000000' y1='1759.000000' x2='5040.000000' y2='1839.000000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='3040.000000' y1='2896.500000' x2='3040.000000' y2='2976.500000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='4840.000000' y1='1040.250000' x2='4840.000000' y2='1120.250000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<line x1='5640.000000' y1='1171.500000' x2='5640.000000' y2='1251.500000' stroke='rgb(51,51,178)' style='stroke-dasharray: 1, 1'  />
<g transform='translate(4489.636364,2159.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>P._afra</text></g>
<g transform='translate(6289.636364,2359.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>P._phoenicoptera</text></g>
<g transform='translate(6689.636364,1059.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._r_cingica</text></g>
<g transform='translate(4689.636364,2959.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._rhodophyga</text></g>
<g transform='translate(1089.636364,59.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>O._atricolis</text></g>
<g transform='translate(1989.636364,359.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>G._granatia</text></g>
<g transform='translate(3289.636364,559.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>H._niveoguttatus</text></g>
<g transform='translate(5889.636364,1559.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._rufopicta</text></g>
<g transform='translate(5289.636364,2259.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>P._lineata</text></g>
<g transform='translate(2689.636364,459.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._dybowskii</text></g>
<g transform='translate(4389.636364,2059.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>P._melba_citerior</text></g>
<g transform='translate(6889.636364,1259.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._virata</text></g>
<g transform='translate(4889.636364,859.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._larvata</text></g>
<g transform='translate(3389.636364,659.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>H._margaritatus</text></g>
<g transform='translate(5589.636364,3159.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._melpoda</text></g>
<g transform='translate(5689.636364,959.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._rara</text></g>
<g transform='translate(4289.636364,1959.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>P._melba_grotei</text></g>
<g transform='translate(3089.636364,2759.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._astrild</text></g>
<g transform='translate(1189.636364,159.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>A._subflava</text></g>
<g transform='translate(2389.636364,2659.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>C._melanotis</text></g>
<g transform='translate(3489.636364,759.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>C._monteiri</text></g>
<g transform='translate(6389.636364,2459.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>P._hypogrammica</text></g>
<g transform='translate(5989.636364,1659.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._nitidula</text></g>
<g transform='translate(2289.636364,2559.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>C._quartinia</text></g>
<g transform='translate(7189.636364,1459.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._sanguinodorsalis</text></g>
<g transform='translate(1889.636364,259.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>G._ianthinogaster</text></g>
<g transform='translate(6189.636364,1859.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._senegala_rhodopsis</text></g>
<g transform='translate(2589.636364,3259.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._erythronotos</text></g>
<g transform='translate(3889.636364,2859.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._paludicola</text></g>
<g transform='translate(6789.636364,1159.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._r._rubricata</text></g>
<g transform='translate(6089.636364,1759.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._senegala_rendalii</text></g>
<g transform='translate(7089.636364,1359.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>L._rhodopareia</text></g>
<g transform='translate(5489.636364,3059.000000) rotate(0.000000)'><text x='0' y='0' font-size='20.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(51,51,178)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>E._troglodytes</text></g>
<line x1='6240.000000' y1='2449.000000' x2='5240.000000' y2='2399.000000' stroke='rgb(0,0,0)'  />
<line x1='7000.000000' y1='1439.000000' x2='6960.000000' y2='1429.000000' stroke='rgb(0,0,0)'  />
<line x1='1840.000000' y1='349.000000' x2='1340.000000' y2='299.000000' stroke='rgb(0,0,0)'  />
<path d='M2890.000000 574.000000 C4878.333333 969.833333 4878.333333 969.833333 6906.666667 1365.666667'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='2440.000000' y1='3249.000000' x2='1640.000000' y2='3045.875000' stroke='rgb(0,0,0)'  />
<path d='M5440.000000 3149.000000 C4020.000000 2972.437500 4020.000000 2972.437500 2640.000000 2795.875000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='1990.000000' y1='2944.312500' x2='1640.000000' y2='3045.875000' stroke='rgb(0,0,0)'  />
<line x1='6906.666667' y1='1365.666667' x2='6873.333333' y2='1382.333333' stroke='rgb(0,0,0)'  />
<path d='M5540.000000 949.000000 C6250.000000 1194.000000 6250.000000 1194.000000 7000.000000 1439.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='1040.000000' y1='149.000000' x2='740.000000' y2='99.000000' stroke='rgb(0,0,0)'  />
<line x1='2340.000000' y1='2842.750000' x2='1990.000000' y2='2944.312500' stroke='rgb(0,0,0)'  />
<line x1='2640.000000' y1='2795.875000' x2='2340.000000' y2='2842.750000' stroke='rgb(0,0,0)'  />
<path d='M3540.000000 1999.000000 C2745.000000 2471.656250 2745.000000 2471.656250 1990.000000 2944.312500'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='6140.000000' y1='2349.000000' x2='5240.000000' y2='2399.000000' stroke='rgb(0,0,0)'  />
<path d='M5240.000000 2399.000000 C4545.000000 2211.500000 4545.000000 2211.500000 3890.000000 2024.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='940.000000' y1='49.000000' x2='740.000000' y2='99.000000' stroke='rgb(0,0,0)'  />
<line x1='1740.000000' y1='249.000000' x2='1340.000000' y2='299.000000' stroke='rgb(0,0,0)'  />
<line x1='6940.000000' y1='1349.000000' x2='6906.666667' y2='1365.666667' stroke='rgb(0,0,0)'  />
<path d='M6040.000000 1849.000000 C6320.000000 1605.250000 6320.000000 1605.250000 6640.000000 1361.500000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='6960.000000' y1='1429.000000' x2='6920.000000' y2='1419.000000' stroke='rgb(0,0,0)'  />
<path d='M6640.000000 1149.000000 C6736.666667 1265.666667 6736.666667 1265.666667 6873.333333 1382.333333'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='2940.000000' y1='2749.000000' x2='2640.000000' y2='2795.875000' stroke='rgb(0,0,0)'  />
<line x1='3140.000000' y1='549.000000' x2='2890.000000' y2='574.000000' stroke='rgb(0,0,0)'  />
<path d='M740.000000 99.000000 C3790.000000 754.000000 3790.000000 754.000000 6880.000000 1409.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <path d='M5940.000000 1749.000000 C4395.000000 1161.500000 4395.000000 1161.500000 2890.000000 574.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='6840.000000' y1='1399.000000' x2='6640.000000' y2='1361.500000' stroke='rgb(0,0,0)'  />
<line x1='6880.000000' y1='1409.000000' x2='6840.000000' y2='1399.000000' stroke='rgb(0,0,0)'  />
<line x1='6873.333333' y1='1382.333333' x2='6840.000000' y2='1399.000000' stroke='rgb(0,0,0)'  />
<line x1='6920.000000' y1='1419.000000' x2='6880.000000' y2='1409.000000' stroke='rgb(0,0,0)'  />
<line x1='3840.000000' y1='1974.000000' x2='3540.000000' y2='1999.000000' stroke='rgb(0,0,0)'  />
<line x1='3890.000000' y1='2024.000000' x2='3540.000000' y2='1999.000000' stroke='rgb(0,0,0)'  />
<line x1='7040.000000' y1='1449.000000' x2='7000.000000' y2='1439.000000' stroke='rgb(0,0,0)'  />
<line x1='4240.000000' y1='2049.000000' x2='3890.000000' y2='2024.000000' stroke='rgb(0,0,0)'  />
<line x1='4140.000000' y1='1949.000000' x2='3840.000000' y2='1974.000000' stroke='rgb(0,0,0)'  />
<line x1='1340.000000' y1='299.000000' x2='1240.000000' y2='487.134766' stroke='rgb(0,0,0)'  />
<path d='M6640.000000 1361.500000 C3920.000000 924.317383 3920.000000 924.317383 1240.000000 487.134766'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <path d='M1240.000000 487.134766 C1320.000000 1710.645508 1320.000000 1710.645508 1440.000000 2934.156250'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <line x1='1640.000000' y1='3045.875000' x2='1440.000000' y2='2934.156250' stroke='rgb(0,0,0)'  />
<path d='M5740.000000 1549.000000 C6310.000000 1484.000000 6310.000000 1484.000000 6920.000000 1419.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <path d='M4340.000000 2149.000000 C4070.000000 2061.500000 4070.000000 2061.500000 3840.000000 1974.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <path d='M3340.000000 749.000000 C5130.000000 1089.000000 5130.000000 1089.000000 6960.000000 1429.000000'  style='stroke-dasharray: 4, 2' stroke='rgb(0,0,0)' fill='rgb(0,0,0)' fill-opacity='0.000000'  />
 <rect x='6995.000000' y='1434.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6995.000000,1434.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='2885.000000' y='569.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(2885.000000,569.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='1985.000000' y='2939.312500' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(1985.000000,2939.312500) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6901.666667' y='1360.666667' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6901.666667,1360.666667) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='2335.000000' y='2837.750000' width='10.000000' height='10.000000' stroke='rgb(127,127,127)' fill='rgb(255,255,255)'  stroke-width='1.000000'/>
<g transform='translate(2335.000000,2837.750000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,255)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='2635.000000' y='2790.875000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(2635.000000,2790.875000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='3535.000000' y='1994.000000' width='10.000000' height='10.000000' stroke='rgb(0,0,0)' fill='rgb(0,0,0)'  stroke-width='1.000000'/>
<g transform='translate(3535.000000,1994.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='5235.000000' y='2394.000000' width='10.000000' height='10.000000' stroke='rgb(0,0,0)' fill='rgb(0,0,0)'  stroke-width='1.000000'/>
<g transform='translate(5235.000000,2394.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6955.000000' y='1424.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6955.000000,1424.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='735.000000' y='94.000000' width='10.000000' height='10.000000' stroke='rgb(0,0,0)' fill='rgb(0,0,0)'  stroke-width='1.000000'/>
<g transform='translate(735.000000,94.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6835.000000' y='1394.000000' width='10.000000' height='10.000000' stroke='rgb(0,0,0)' fill='rgb(0,0,0)'  stroke-width='1.000000'/>
<g transform='translate(6835.000000,1394.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6875.000000' y='1404.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6875.000000,1404.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6868.333333' y='1377.333333' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6868.333333,1377.333333) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6915.000000' y='1414.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6915.000000,1414.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='3835.000000' y='1969.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(3835.000000,1969.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='3885.000000' y='2019.000000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(3885.000000,2019.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='1435.000000' y='2929.156250' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(1435.000000,2929.156250) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='1335.000000' y='294.000000' width='10.000000' height='10.000000' stroke='rgb(0,0,0)' fill='rgb(0,0,0)'  stroke-width='1.000000'/>
<g transform='translate(1335.000000,294.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='6635.000000' y='1356.500000' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(6635.000000,1356.500000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='1235.000000' y='482.134766' width='10.000000' height='10.000000' stroke='rgb(127,127,0)' fill='rgb(255,255,0)'  stroke-width='1.000000'/>
<g transform='translate(1235.000000,482.134766) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(255,255,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<rect x='1635.000000' y='3040.875000' width='10.000000' height='10.000000' stroke='rgb(0,0,0)' fill='rgb(0,0,0)'  stroke-width='1.000000'/>
<g transform='translate(1635.000000,3040.875000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>1.0</text></g>
<g transform='translate(6250.000000,2455.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._togoensis</text></g>
<g transform='translate(1850.000000,355.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._regia</text></g>
<g transform='translate(2450.000000,3255.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._hypocherina</text></g>
<g transform='translate(5450.000000,3155.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._macroura_W.</text></g>
<g transform='translate(5550.000000,955.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._camerunensis</text></g>
<g transform='translate(1050.000000,155.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._raricola</text></g>
<g transform='translate(6150.000000,2355.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._interjecta</text></g>
<g transform='translate(950.000000,55.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._nigeriae</text></g>
<g transform='translate(1750.000000,255.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._fischeri</text></g>
<g transform='translate(6950.000000,1355.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._purpurascens</text></g>
<g transform='translate(6050.000000,1855.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._chalybeata_W.</text></g>
<g transform='translate(6650.000000,1155.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._funera</text></g>
<g transform='translate(2950.000000,2755.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._macroura_S</text></g>
<g transform='translate(3150.000000,555.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._codringtoni</text></g>
<g transform='translate(5950.000000,1755.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._chalybeata_S.</text></g>
<g transform='translate(7050.000000,1455.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._maryae</text></g>
<g transform='translate(4250.000000,2055.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._orientalis</text></g>
<g transform='translate(4150.000000,1955.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._paradisaea</text></g>
<g transform='translate(5750.000000,1555.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._wilsoni</text></g>
<g transform='translate(4350.000000,2155.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._obtusa</text></g>
<g transform='translate(3350.000000,755.000000) rotate(0.000000)'><text x='0' y='0' font-size='14.000000' stroke='rgb(0,0,0)' stroke-opacity='0.000000' fill='rgb(0,0,0)'  stroke-width='1.000000' text-anchor='start' style='dominant-baseline: auto'>V._larvaticola</text></g>
</g>
</g>
</g></svg>